----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:37:02 05/15/2018 
-- Design Name: 
-- Module Name:    DAC_8_bit - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity DAC_8_bit is
    Port ( i_clk : in  STD_LOGIC;
           in_rst : in  STD_LOGIC;
			  i_slv_4: in std_logic_vector( 31 downto 0);
           o_strobe : out  STD_LOGIC;
           o_clk : out  STD_LOGIC;
           o_data : out  STD_LOGIC_vector (7 downto 0));
end DAC_8_bit;

architecture Behavioral of DAC_8_bit is

begin


end Behavioral;

